library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.NUMERIC_STD.ALL; 

entity RAM is
port(
    clk         : in  std_logic; 
    Adress      : in  std_logic_vector(7 downto 0);
    Data_in     : in  std_logic_vector(23 downto 0);
    EnRAM       : in  std_logic; 
    RW          : in  std_logic; 
    j1, j2      : in  STD_LOGIC_VECTOR(0 to 8);
    gana        : in  std_logic_vector(1 downto 0);
    ganador, empat, ini : in std_logic;
    sumar2      : in  std_logic_vector(1 downto 0);
    torneo      : in  std_logic;
    Data_out    : out std_logic_vector(23 downto 0)
);
end RAM;

architecture Behavioral of RAM is
    signal sum2: std_logic_vector(1 downto 0);
    signal col0_dyn, col3_dyn, col6_dyn : std_logic_vector(7 downto 0);
    signal status_byte : std_logic_vector(7 downto 0);
    signal addr_int : integer range 0 to 255; 

    type RAM_MEMORY is array (0 to 255) of std_logic_vector(23 downto 0);
    
    signal MEMORY: RAM_MEMORY := (
        -- 1. MENU
        0 => "00001011" & "00000001" & "11010110", 
        1 => "00011111" & "00000001" & "00010100", 
        2 => "00010010" & "00000000" & "00001010", 
        
        -- MODO TORNEO
        3 => "00001011" & "00001000" & "11001010", 
        4 => "00001011" & "00001001" & "11001010", 
        5 => "00001011" & "00001010" & "11001010", 
        6 => "00001011" & "00001011" & "11001010", 
        7 => "00001011" & "00001100" & "11001010", 
        8 => "00001011" & "00001101" & "11001010", 
        9 => "00001011" & "00001110" & "11001010", 
        10=> "00001011" & "00001111" & "11001010", 
        11=> "00000001" & "00000101" & "00000101", 
        12=> "00010000" & "00000000" & "00000000", 

        -- MODO NORMAL
        13 => "00011111" & "00000001" & "00000100", 
        14 => "00010010" & "00000000" & "00001010", 
        15 => "00001011" & "00001000" & "11101000", 
        16 => "00001011" & "00001001" & "11101000", 
        17 => "00001011" & "00001010" & "11101000", 
        18 => "00001011" & "00001011" & "11101000", 
        19 => "00001011" & "00001100" & "11101000", 
        20 => "00001011" & "00001101" & "11101000", 
        21 => "00001011" & "00001110" & "11101000", 
        22 => "00001011" & "00001111" & "11101000", 
        23=> "00000001" & "00000101" & "00000101", 
        24=> "00010000" & "00000000" & "00000000", 

        -- 2. JUEGO
        -- Empate
        25=> "00011111" & "00000001" & "00000010", 
        26=> "00010010" & "00000000" & "00001011", 
        27=> "00001011" & "00001000" & "10111100", 
        28=> "00001011" & "00001001" & "10111100", 
        29=> "00001011" & "00001010" & "10111100", 
        30=> "00001011" & "00001011" & "10111100", 
        31=> "00001011" & "00001100" & "10111100", 
        32=> "00001011" & "00001101" & "10111100", 
        33=> "00001011" & "00001110" & "10111100", 
        34=> "00001011" & "00001111" & "10111100", 
        35=> "00000001" & "00000101" & "00000101", 
        36=> "00010000" & "00000000" & "00000000", 
        37=> "00011010" & "00000000" & "00000000", 

        -- Ganador J1
        38=> "00011111" & "00000001" & "00000001", 
        39=> "00010010" & "00000000" & "00001101", 
        40=> "00011111" & "00000101" & "00000001", 
        41=> "00010011" & "00000000" & "00000010", 
        42=> "00011011" & "00000110" & "00001010", 
        43=> "00011011" & "00000101" & "00000001", 
        44=> "00001011" & "00001000" & "10111011", 
        45=> "00001011" & "00001001" & "10111011", 
        46=> "00001011" & "00001010" & "10111011", 
        47=> "00001011" & "00001011" & "10111011", 
        48=> "00001011" & "00001100" & "10111011", 
        49=> "00001011" & "00001101" & "10111011", 
        50=> "00001011" & "00001110" & "10111011", 
        51=> "00001011" & "00001111" & "10111011", 
        52=> "00010000" & "00000000" & "00000000", 

        -- Ganador J2
        53=> "00011111" & "00000001" & "00001001", 
        54=> "00010010" & "00000000" & "00001101", 
        55=> "00011111" & "00000101" & "00000001", 
        56=> "00010011" & "00000000" & "00000010", 
        57=> "00011011" & "00000111" & "00001010", 
        58=> "00011011" & "00000101" & "00000001", 
        59=> "00001011" & "00001000" & "10100100", 
        60=> "00001011" & "00001001" & "10100100", 
        61=> "00001011" & "00001010" & "10100100", 
        62=> "00001011" & "00001011" & "10100100", 
        63=> "00001011" & "00001100" & "10100100", 
        64=> "00001011" & "00001101" & "10100100", 
        65=> "00001011" & "00001110" & "10100100", 
        66=> "00001011" & "00001111" & "10100100", 
        67=> "00010000" & "00000000" & "00000000", 

        -- Default
        68=> "00000001" & "00000101" & "00000101", 
        69=> "00001011" & "00001000" & "10101010", 
        70=> "00001011" & "00001001" & "10101010", 
        71=> "00001011" & "00001010" & "10101010", 
        72=> "00001011" & "00001011" & "10101010", 
        73=> "00001011" & "00001100" & "10101010", 
        74=> "00001011" & "00001101" & "10101010", 
        75=> "00001011" & "00001110" & "10101010", 
        76=> "00001011" & "00001111" & "10101010", 
        
        -- Suma Movimiento
        77=> "00001011" & "00000100" & "10001000", 
        78=> "00011111" & "00000100" & "00000000", 
        79=> "00010010" & "00000000" & "00000011", 
        80=> "00000001" & "00000011" & "00000011", 
        81=> "00010000" & "00000000" & "00000000", 
        82=> "00011010" & "00000000" & "00000000", 

        -- Check Fin Torneo (3)
        83=> "00011111" & "00000100" & "00000011", 
        84=> "00010010" & "00000000" & "00000010", -- BNZ 87
        
        -- CORREGIDO: JMP 130 (10000010)
        85=> "00010000" & "00000000" & "10000010", -- JMP 130
        86=> "00011010" & "00000000" & "00000000", 

        -- J1 Move
        87=> "00011111" & "00000100" & "00000001", 
        88=> "00010010" & "00000000" & "00000101", 
        89=> "00011111" & "00000011" & "00000001",
        90=> "00010011" & "00000000" & "00001000",
        91=> "00011011" & "00000110" & "00000010", 
        92=> "00011011" & "00000011" & "00000001",
        93=> "00010000" & "00000000" & "00000000", 
        
        -- J2 Move
        94=> "00011111" & "00000011" & "00000001",
        95=> "00010011" & "00000000" & "00000011",
        96=> "00011011" & "00000111" & "00000010",
        97=> "00011011" & "00000011" & "00000001",
        98=> "00010000" & "00000000" & "00000000", 
        99=> "00010000" & "00000000" & "00000000", 

        -- CEREMONIA (130)
        130=> "00000100" & "00000110" & "00000111", -- CMP R6, R7
        131=> "00010100" & "00000000" & "00001001", -- BS1 -> 141
        
        -- Gana J1
        132=> "00001011" & "00001000" & "00011100", -- LW R8, [160]
        133=> "00001011" & "00001001" & "00011100", 
        134=> "00001011" & "00001010" & "00011100", 
        135=> "00001011" & "00001011" & "00011100", 
        136=> "00001011" & "00001100" & "00011100", 
        137=> "00001011" & "00001101" & "00011100", 
        138=> "00001011" & "00001110" & "00011100", 
        139=> "00001011" & "00001111" & "00011100", 
        140=> "00010000" & "00000000" & "10000010", -- Loop 130

        -- Gana J2
        141=> "00001011" & "00001000" & "00010111", -- LW R8, [168]
        142=> "00001011" & "00001001" & "00010111", 
        143=> "00001011" & "00001010" & "00010111", 
        144=> "00001011" & "00001011" & "00010111", 
        145=> "00001011" & "00001100" & "00010111", 
        146=> "00001011" & "00001101" & "00010111", 
        147=> "00001011" & "00001110" & "00010111", 
        148=> "00001011" & "00001111" & "00010111", 
        149=> "00010000" & "00000000" & "10001101", -- Loop 141

        -- DATOS
        -- J1 (160: Apagado)
        160 => "00000000" & "00000000" & "00000000",
        161 => "00000000" & "00000000" & "00000000",
        162 => "00000000" & "00000000" & "00000000",
        163 => "00000000" & "00000000" & "00000000",
        164 => "00000000" & "00000000" & "00000000",
        165 => "00000000" & "00000000" & "00000000",
        166 => "00000000" & "00000000" & "00000000",
        167 => "00000000" & "00000000" & "00000000",

        -- J2 (168: Encendido)
        168 => "00000000" & "00000000" & "11111111",
        169 => "00000000" & "00000000" & "11111111",
        170 => "00000000" & "00000000" & "11111111",
        171 => "00000000" & "00000000" & "11111111",
        172 => "00000000" & "00000000" & "11111111",
        173 => "00000000" & "00000000" & "11111111",
        174 => "00000000" & "00000000" & "11111111",
        175 => "00000000" & "00000000" & "11111111",

        -- (Resto de Datos: 206 en adelante IGUAL QUE ANTES)
        206 => "00000000" & "00000000" & "10000111",
        -- ... (Manten el resto de tus datos aqui) ...
        
        -- Para que no se te pierdan los datos si copias:
        207 => "00000000" & "00000000" & "01111011",
        208 => "00000000" & "00000000" & "10000010",
        209 => "00000000" & "00000000" & "11000000",
        210 => "00000000" & "00000000" & "11000000",
        211 => "00000000" & "00000000" & "10000010",
        212 => "00000000" & "00000000" & "01111011",
        213 => "00000000" & "00000000" & "10000111",
        
        216 => "00000000" & "00000000" & "00000000",
        217 => "00000000" & "00000000" & "01111110",
        218 => "00000000" & "00000000" & "01011010",
        219 => "00000000" & "00000000" & "01011010",
        220 => "00000000" & "00000000" & "01011010",
        221 => "00000000" & "00000000" & "01011010",
        222 => "00000000" & "00000000" & "01111110",
        223 => "00000000" & "00000000" & "00000000",

        224 => "00000000" & "00000000" & "00000000",
        225 => "00000000" & "00000000" & "01111110",
        226 => "00000000" & "00000000" & "01111010",
        227 => "00000000" & "00000000" & "01010010",
        228 => "00000000" & "00000000" & "01111110",
        229 => "00000000" & "00000000" & "01010010",
        230 => "00000000" & "00000000" & "01001010",
        231 => "00000000" & "00000000" & "00000000",

        232 => "00000000" & "00000000" & "00000000",
        233 => "00000000" & "00000000" & "01111110",
        234 => "00000000" & "00000000" & "01111010",
        235 => "00000000" & "00000000" & "01010010",
        236 => "00000000" & "00000000" & "01111110",
        237 => "00000000" & "00000000" & "01000010",
        238 => "00000000" & "00000000" & "01111110",
        239 => "00000000" & "00000000" & "00000000",

        240 => "00000000" & "00000000" & "11011011",
        241 => "00000000" & "00000000" & "11011011",
        242 => "00000000" & "00000000" & "00000000",
        243 => "00000000" & "00000000" & "11011011",
        244 => "00000000" & "00000000" & "11011011",
        245 => "00000000" & "00000000" & "00000000",
        246 => "00000000" & "00000000" & "11011011",
        247 => "00000000" & "00000000" & "11011011",

        248 => "00000000" & "00000000" & "00011110",
        249 => "00000000" & "00000000" & "10101001",
        250 => "00000000" & "00000000" & "10010000",
        251 => "00000000" & "00000000" & "10101000",
        252 => "00000000" & "00000000" & "00011000",
        253 => "00000000" & "00000000" & "11111100",
        254 => "00000000" & "00000000" & "11111110",
        255 => "00000000" & "00000000" & "11000001",

        others => (others => '0')
    );
 
begin
    addr_int <= to_integer(unsigned(Adress));
    sum2<=sumar2;

    col0_dyn <= j1(0) & j2(0) & '0' & j1(3) & j2(3) & '0' & j1(6) & j2(6);
    col3_dyn <= j1(1) & j2(1) & '0' & j1(4) & j2(4) & '0' & j1(7) & j2(7);
    col6_dyn <= j1(2) & j2(2) & '0' & j1(5) & j2(5) & '0' & j1(8) & j2(8);

    status_byte <= "000" & (torneo and ini) & gana(1) & ini & empat & ganador;

    process(addr_int, MEMORY, col0_dyn, col3_dyn, col6_dyn, status_byte, sum2)
    begin
        case addr_int is
            when 214 => Data_out <= x"0000" & "000000"&sum2; 
            when 215 => Data_out <= x"0000" & status_byte;
            when 240 => Data_out <= x"0000" & col0_dyn;
            when 243 => Data_out <= x"0000" & col3_dyn;
            when 246 => Data_out <= x"0000" & col6_dyn;
            when others => Data_out <= MEMORY(addr_int);
        end case;
    end process;

    process(clk)
    begin
        if rising_edge(clk) then
            if EnRAM = '1' and RW = '0' then 
                MEMORY(addr_int) <= Data_in;
            end if;
        end if;
    end process;

end Behavioral;