library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.NUMERIC_STD.ALL; 

entity RAM is
port(
    clk         : in  std_logic; 
    Adress      : in  std_logic_vector(7 downto 0);
    Data_in     : in  std_logic_vector(23 downto 0);
    EnRAM       : in  std_logic; 
    RW          : in  std_logic; 
    j1, j2      : in  STD_LOGIC_VECTOR(0 to 8);
    gana        : in  std_logic_vector(1 downto 0);
    ganador, empat, ini : in std_logic;
    sumar2      : in  std_logic_vector(1 downto 0);
    torneo      : in  std_logic;
    Data_out    : out std_logic_vector(23 downto 0)
);
end RAM;

architecture Behavioral of RAM is
    signal sum2: std_logic_vector(1 downto 0);
    signal col0_dyn, col3_dyn, col6_dyn : std_logic_vector(7 downto 0);
    signal status_byte : std_logic_vector(7 downto 0);
    signal addr_int : integer range 0 to 255; 

    type RAM_MEMORY is array (0 to 255) of std_logic_vector(23 downto 0);
    
    signal MEMORY: RAM_MEMORY := (
        -- ==========================================================
        -- 1. MENU (Check 80)
        -- ==========================================================
        0 => "00001011" & "00000001" & "11010110", -- LW R1, [Estado]
        1 => "00011111" & "00000001" & "01010000", -- CMPI R1, 80
        2 => "00010010" & "00000000" & "00001010", -- BNZ 13 (A Modo Normal)
        
        -- Carga Imagen Torneo (Menu)
        3 => "00001011" & "00001000" & "11001010", -- LW R8
        4 => "00001011" & "00001001" & "11001010", 
        5 => "00001011" & "00001010" & "11001010", 
        6 => "00001011" & "00001011" & "11001010", 
        7 => "00001011" & "00001100" & "11001010", 
        8 => "00001011" & "00001101" & "11001010", 
        9 => "00001011" & "00001110" & "11001010", 
        10=> "00001011" & "00001111" & "11001010", 
        11=> "00000001" & "00000101" & "00000101", -- Reset Flags
        12=> "00010000" & "00000000" & "00000000", -- JMP 0

        -- ==========================================================
        -- 2. MODO NORMAL (Check 16)
        -- ==========================================================
        13 => "00011111" & "00000001" & "00010000", -- CMPI R1, 16
        14 => "00010010" & "00000000" & "00001010", -- BNZ 25 (A Empate)
        
        -- Carga Imagen Normal Inicial
        15 => "00001011" & "00001000" & "11101000", -- LW R8
        16 => "00001011" & "00001001" & "11101000", 
        17 => "00001011" & "00001010" & "11101000", 
        18 => "00001011" & "00001011" & "11101000", 
        19 => "00001011" & "00001100" & "11101000", 
        20 => "00001011" & "00001101" & "11101000", 
        21 => "00001011" & "00001110" & "11101000", 
        22 => "00001011" & "00001111" & "11101000", 
        23=> "00000001" & "00000101" & "00000101", 
        24=> "00010000" & "00000000" & "00000000", -- JMP 0

        -- ==========================================================
        -- 3. CHECK EMPATE (Check 8)
        -- ==========================================================
        25=> "00011111" & "00000001" & "00001000", -- CMPI R1, 8
        26=> "00010010" & "00000000" & "00001011", -- BNZ 38 (A Check Fin Torneo)
        
        -- Carga Imagen Empate
        27=> "00001011" & "00001000" & "10111100", 
        28=> "00001011" & "00001001" & "10111100", 
        29=> "00001011" & "00001010" & "10111100", 
        30=> "00001011" & "00001011" & "10111100", 
        31=> "00001011" & "00001100" & "10111100", 
        32=> "00001011" & "00001101" & "10111100", 
        33=> "00001011" & "00001110" & "10111100", 
        34=> "00001011" & "00001111" & "10111100", 
        35=> "00000001" & "00000101" & "00000101", 
        36=> "00010000" & "00000000" & "00000000", -- JMP 0
        37=> "00011010" & "00000000" & "00000000", -- NOP

        -- ==========================================================
        -- 4. CHECK FIN TORNEO UNIVERSAL (Lines 38-60)
        -- ==========================================================
        -- Cargamos sumar2 desde la dirección 214
        -- Offset: 214 - 39 = 175 = 10101111
        38=> "00001011" & "00000100" & "10101111", -- LW R4, [214]
        
        -- Verificamos si es 3 (Fin de Torneo)
        39=> "00011111" & "00000100" & "00000011", -- CMPI R4, 3
        
        -- Si NO es 3, saltamos a la lógica normal (J1 Normal)
        -- Offset: 61 - 41 = 20 = 00010100
        40=> "00010010" & "00000000" & "00010100", -- BNZ 61 (A J1 Normal)

        -- === SÍ ES FIN DE TORNEO (Ganador o Empate) ===
        -- Comparamos puntajes (R6 vs R7)
        41=> "00000100" & "00000110" & "00000111", -- CMP R6, R7
        
        -- Si R6 < R7 (J2 gana), saltamos a cargar J2
        -- Offset: 52 - 43 = 9 = 00001001
        42=> "00010100" & "00000000" & "00001001", -- BS1 52 (A J2 Torneo)

        -- GANA J1 TORNEO (Cargar 160)
        -- Offset: 160 - 44 = 116 = 01110100
        43=> "00001011" & "00001000" & "01110100", -- LW R8, [160]
        44=> "00001011" & "00001001" & "01110100", 
        45=> "00001011" & "00001010" & "01110100", 
        46=> "00001011" & "00001011" & "01110100", 
        47=> "00001011" & "00001100" & "01110100", 
        48=> "00001011" & "00001101" & "01110100", 
        49=> "00001011" & "00001110" & "01110100", 
        50=> "00001011" & "00001111" & "01110100", 
        51=> "00100100" & "00000000" & "00000000", -- HALT J1

        -- GANA J2 TORNEO (Cargar 168)
        -- Offset: 168 - 53 = 115 = 01110011
        52=> "00001011" & "00001000" & "01110011", -- LW R8, [168]
        53=> "00001011" & "00001001" & "01110011", 
        54=> "00001011" & "00001010" & "01110011", 
        55=> "00001011" & "00001011" & "01110011", 
        56=> "00001011" & "00001100" & "01110011", 
        57=> "00001011" & "00001101" & "01110011", 
        58=> "00001011" & "00001110" & "01110011", 
        59=> "00001011" & "00001111" & "01110011", 
        60=> "00100100" & "00000000" & "00000000", -- HALT J2

        -- ==========================================================
        -- 5. CHECK GANADOR J1 NORMAL (Check 4)
        -- ==========================================================
        61=> "00011111" & "00000001" & "00000100", -- CMPI R1, 4
        62=> "00010010" & "00000000" & "00001101", -- BNZ 76 (A J2 Normal)
        
        -- Suma Puntos
        63=> "00011111" & "00000101" & "00000001", -- CMPI R5, 1
        64=> "00010011" & "00000000" & "00000010", -- BZ +2
        65=> "00011011" & "00000110" & "00001010", -- ADDI R6, 10
        66=> "00011011" & "00000101" & "00000001", -- ADDI R5, 1
        
        -- Carga J1 Normal (232)
        -- Offset: 232 - 68 = 164 = 10100100
        67=> "00001011" & "00001000" & "10100100", -- LW R8, [232]
        68=> "00001011" & "00001001" & "10100100", 
        69=> "00001011" & "00001010" & "10100100", 
        70=> "00001011" & "00001011" & "10100100", 
        71=> "00001011" & "00001100" & "10100100", 
        72=> "00001011" & "00001101" & "10100100", 
        73=> "00001011" & "00001110" & "10100100", 
        74=> "00001011" & "00001111" & "10100100", 
        75=> "00010000" & "00000000" & "00000000", -- JMP 0

        -- ==========================================================
        -- 6. CHECK GANADOR J2 NORMAL (Check 36)
        -- ==========================================================
        76=> "00011111" & "00000001" & "00100100", -- CMPI R1, 36
        77=> "00010010" & "00000000" & "00001101", -- BNZ 91 (A Default)
        
        -- Suma Puntos
        78=> "00011111" & "00000101" & "00000001", 
        79=> "00010011" & "00000000" & "00000010", 
        80=> "00011011" & "00000111" & "00001010", 
        81=> "00011011" & "00000101" & "00000001", 
        
        -- Carga J2 Normal (224)
        -- Offset: 224 - 83 = 141 = 10001101
        82=> "00001011" & "00001000" & "10001101", -- LW R8, [224]
        83=> "00001011" & "00001001" & "10001101", 
        84=> "00001011" & "00001010" & "10001101", 
        85=> "00001011" & "00001011" & "10001101", 
        86=> "00001011" & "00001100" & "10001101", 
        87=> "00001011" & "00001101" & "10001101", 
        88=> "00001011" & "00001110" & "10001101", 
        89=> "00001011" & "00001111" & "10001101", 
        90=> "00010000" & "00000000" & "00000000", -- JMP 0

        -- ==========================================================
        -- 7. DEFAULT / JUEGO EN CURSO
        -- ==========================================================
        91=> "00000001" & "00000101" & "00000101", -- SUB R5, R5
        
        -- LOAD TABLERO (240)
        -- Offset: 240 - 93 = 147 = 10010011
        92=> "00001011" & "00001000" & "10010011", -- LW R8
        93=> "00001011" & "00001001" & "10010011", 
        94=> "00001011" & "00001010" & "10010011", 
        95=> "00001011" & "00001011" & "10010011", 
        96=> "00001011" & "00001100" & "10010011", 
        97=> "00001011" & "00001101" & "10010011", 
        98=> "00001011" & "00001110" & "10010011", 
        99=> "00001011" & "00001111" & "10010011", 
        
        -- SUMA MOV (Desde 100)
        100=> "00001011" & "00000100" & "01110001", -- LW R4, [214] (Offset: 214-101=113)
        101=> "00011111" & "00000100" & "00000000", -- CMPI R4, 0
        102=> "00010010" & "00000000" & "00000011", -- BNZ 106
        103=> "00000001" & "00000011" & "00000011", -- SUB R3, R3
        104=> "00010000" & "00000000" & "00000000", -- JMP 0
        105=> "00011010" & "00000000" & "00000000", -- NOP

        -- MOV J1
        106=> "00011111" & "00000100" & "00000001", -- CMPI R4, 1
        107=> "00010010" & "00000000" & "00000101", -- BNZ 113
        108=> "00011111" & "00000011" & "00000001", -- CMPI R3, 1
        109=> "00010011" & "00000000" & "00001000", -- BZ 118
        110=> "00011011" & "00000110" & "00000010", -- ADDI R6, 2
        111=> "00011011" & "00000011" & "00000001", -- ADDI R3, 1
        112=> "00010000" & "00000000" & "00000000", -- JMP 0
        
        -- MOV J2
        113=> "00011111" & "00000011" & "00000001", -- CMPI R3, 1
        114=> "00010011" & "00000000" & "00000011", -- BZ 118
        115=> "00011011" & "00000111" & "00000010", -- ADDI R7, 2
        116=> "00011011" & "00000011" & "00000001", -- ADDI R3, 1
        117=> "00010000" & "00000000" & "00000000", -- JMP 0
        118=> "00010000" & "00000000" & "00000000", -- JMP 0

        -- ==========================================================
        -- DATOS Y PATRONES
        -- ==========================================================
        
       -- 160-167: J1 GANA TORNEO
        160 => "00000000" & "00000000" & "11000011", 
        161 => "00000000" & "00000000" & "10111101",
        162 => "00000000" & "00000000" & "01111110",
        163 => "00000000" & "00000000" & "01011110",
        164 => "00000000" & "00000000" & "01000010",
        165 => "00000000" & "00000000" & "01111110",
        166 => "00000000" & "00000000" & "10111101",
        167 => "00000000" & "00000000" & "11000011",

        -- 168-175: J2 GANA TORNEO
        168 => "00000000" & "00000000" & "11000011",
        169 => "00000000" & "00000000" & "10111101",
        170 => "00000000" & "00000000" & "01111110",
        171 => "00000000" & "00000000" & "01010010",
        172 => "00000000" & "00000000" & "01001010",
        173 => "00000000" & "00000000" & "01111110",
        174 => "00000000" & "00000000" & "10111101",
        175 => "00000000" & "00000000" & "11000011",
        -- 206 TROFEO
        206 => "00000000" & "00000000" & "10000111",
        207 => "00000000" & "00000000" & "01111011",
        208 => "00000000" & "00000000" & "10000010",
        209 => "00000000" & "00000000" & "11000000",
        210 => "00000000" & "00000000" & "11000000",
        211 => "00000000" & "00000000" & "10000010",
        212 => "00000000" & "00000000" & "01111011",
        213 => "00000000" & "00000000" & "10000111",
        
        -- DATOS EXTRA
        216 => "00000000" & "00000000" & "00000000",
        217 => "00000000" & "00000000" & "01111110",
        218 => "00000000" & "00000000" & "01011010",
        219 => "00000000" & "00000000" & "01011010",
        220 => "00000000" & "00000000" & "01011010",
        221 => "00000000" & "00000000" & "01011010",
        222 => "00000000" & "00000000" & "01111110",
        223 => "00000000" & "00000000" & "00000000",

        -- 224-231 J2 Normal
        224 => "00000000" & "00000000" & "00000000",
        225 => "00000000" & "00000000" & "01111110",
        226 => "00000000" & "00000000" & "01111010",
        227 => "00000000" & "00000000" & "01010010",
        228 => "00000000" & "00000000" & "01111110",
        229 => "00000000" & "00000000" & "01010010",
        230 => "00000000" & "00000000" & "01001010",
        231 => "00000000" & "00000000" & "00000000",

        -- 232-239 J1 Normal
        232 => "00000000" & "00000000" & "00000000",
        233 => "00000000" & "00000000" & "01111110",
        234 => "00000000" & "00000000" & "01111010",
        235 => "00000000" & "00000000" & "01010010",
        236 => "00000000" & "00000000" & "01111110",
        237 => "00000000" & "00000000" & "01000010",
        238 => "00000000" & "00000000" & "01111110",
        239 => "00000000" & "00000000" & "00000000",

        -- TABLERO
        240 => "00000000" & "00000000" & "11011011",
        241 => "00000000" & "00000000" & "11011011",
        242 => "00000000" & "00000000" & "00000000",
        243 => "00000000" & "00000000" & "11011011",
        244 => "00000000" & "00000000" & "11011011",
        245 => "00000000" & "00000000" & "00000000",
        246 => "00000000" & "00000000" & "11011011",
        247 => "00000000" & "00000000" & "11011011",

        -- GATO
        248 => "00000000" & "00000000" & "00011110",
        249 => "00000000" & "00000000" & "10101001",
        250 => "00000000" & "00000000" & "10010000",
        251 => "00000000" & "00000000" & "10101000",
        252 => "00000000" & "00000000" & "00011000",
        253 => "00000000" & "00000000" & "11111100",
        254 => "00000000" & "00000000" & "11111110",
        255 => "00000000" & "00000000" & "11000001",

        others => (others => '0')
    );
 
begin
    addr_int <= to_integer(unsigned(Adress));
    sum2<=sumar2;

    col0_dyn <= j1(0) & j2(0) & '0' & j1(3) & j2(3) & '0' & j1(6) & j2(6);
    col3_dyn <= j1(1) & j2(1) & '0' & j1(4) & j2(4) & '0' & j1(7) & j2(7);
    col6_dyn <= j1(2) & j2(2) & '0' & j1(5) & j2(5) & '0' & j1(8) & j2(8);

    -- CONCATENACIÓN CLAVE
    status_byte <= "0" & (torneo and ini) & gana(1) & ini & empat & ganador & sum2;

    process(addr_int, MEMORY, col0_dyn, col3_dyn, col6_dyn, status_byte, sum2)
    begin
        case addr_int is
            when 214 => Data_out <= x"0000" & "000000"&sum2; 
            when 215 => Data_out <= x"0000" & status_byte;
            when 240 => Data_out <= x"0000" & col0_dyn;
            when 243 => Data_out <= x"0000" & col3_dyn;
            when 246 => Data_out <= x"0000" & col6_dyn;
            when others => Data_out <= MEMORY(addr_int);
        end case;
    end process;

    process(clk)
    begin
        if rising_edge(clk) then
            if EnRAM = '1' and RW = '0' then 
                MEMORY(addr_int) <= Data_in;
            end if;
        end if;
    end process;

end Behavioral;
